// G-pixel info ROM
// 480 * 640
module G_rom
   (
      input wire clk,
      input wire [9:0] pix_x, pix_y,
      output wire G
    );
    
    // Internal signal
    reg [0:154] data;
    reg [9:0] pix_y_reg,pix_x_reg;
    
    always@(posedge clk)
       begin
           pix_x_reg <= pix_x;
           pix_y_reg <= pix_y;
       end
       
    
    
    always@*
       case (pix_y_reg[9:2])
        
	8'h000: data =160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h001: data =160'b1111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h002: data =160'b1111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h003: data =160'b1111111111111111111001111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h004: data =160'b1111111111111111110001111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h005: data =160'b1111111111111111111001111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h006: data =160'b1111111111111111111001111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h007: data =160'b1111111000001111111000111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h008: data =160'b1111101111111011111100111111111111110111111111111111111111111111111111111111111111111111111111111111111001111110000011111111111111111111111111111111111111111111;
8'h009: data =160'b1110111111111111111100011111111111110111111111111111111111111111111111100111111110011111111111111111101111111111111110111111111111111111111111111111111111111111;
8'h00a: data =160'b1101111111111110111110011111111111111011111111111111111111111111111101111111111111111001111111111111111111111111111111101111111111111111111111111111111111111111;
8'h00b: data =160'b1101111111111111011110001111111111111011111111111111111111111111110111111111111111111111011111111101111111111111111111111011111111100000000000000000000000000001;
8'h00c: data =160'b1100111111111111101111001111111111111101111111111111111111111111011111111110000001111111110111111011111111111110111111111101111111000000000000000000000000000001;
8'h00d: data =160'b1100011111111111101111000111111111111111111111111111111111111110111111110000000000001111111011111111111111100000000011111111111111011111111111111111111111111101;
8'h00e: data =160'b1110011111111111110111100011111111111110111111111111111111111011111111100001111100000011111100011111111110000001100000111110111111001111111100110110111111111101;
8'h00f: data =160'b1110001111111111111011100011111111111110111111111111111111110111111110001111111111100011111111111111111100011111111110011111011111001111100111110111010011111101;
8'h010: data =160'b1111000111111111111111110000111111111111011111111111111111100111111100111111111111110001111111111111111101111111111111101111011111001110011110110110111100111101;
8'h011: data =160'b1111100011111111111101110000011111111111111111111111111111001111111001111111111111111001111111111111111001111111111111110111101111001001111111010101111110001101;
8'h012: data =160'b1111100001111111111111011111111111111111101111111111111111001111110111111111111111111001111111111111111011111111111111110111101111010001111111110011001011001101;
8'h013: data =160'b1111110000111111111111111111111111111011111111111111111110001111110111111111111111111101111111111111110111111111111111111011101111010011111111110111101011100101;
8'h014: data =160'b1111111000011111111111111111111111101111111111111111111110011111101111111111111111111101111111111111110111111111111111111111111111010011111111100111011111100101;
8'h015: data =160'b1111111100001111111111111111111111111111111111111111111110011111011111111111110001111110111111111111110111111111100011111101110111011001111111010010010111001101;
8'h016: data =160'b1111111110000111111111111111111101111111111111110111111100011111111111111111111100011110111111111111101111111111110001111101110111001000111110110101111110011101;
8'h017: data =160'b1111111110000011111111111111111111111111111111110111111100111110111111111111111100001110111111111111101111111111111000111101110111001110001110110110101000111101;
8'h018: data =160'b1111111111000000111111111111111111111111111111110111111100111110111111111111111100000111111111111111101111111111110000011101110111001111100001110111000011111101;
8'h019: data =160'b1111111111100000011111111111110111111111110000000111111100111111111111111101111000000111011111111111101111111011100011011101110111001111111111110111111111111101;
8'h01a: data =160'b1111111111110000001111111111110001111110000000000111111000111101111111111100000000110111011111111111111111111000000011011101110111001111111111111111111111111101;
8'h01b: data =160'b1111111111111000000111111111111000000000000000001111111000111101111111111100000000110111011111111111111111111000000011011111110111000000000000000000000000000001;
8'h01c: data =160'b1111111111111100000011111111111000000000000000011111111001111101111111111101111011101111011111111111011111111101111110111111110111111111111111000111111111111111;
8'h01d: data =160'b1111111111111110000000111111111000000000000000001111110000111101111111111110111111001111011111111111011111111110011001111111110011111111111111000111111111111111;
8'h01e: data =160'b1111111111111111000000000000000000000000000000001111100000111111111111111111001110111111011111111111101111111111101111111011111001111111111111000111111111111111;
8'h01f: data =160'b1111111111111111100000000000000000000000000000000111000000011111111111111111110011111101111111111111110011111111111111110111111110111111111111000111111111111111;
8'h020: data =160'b1111111111111111110000000000000000000000000000000010011111111101111111111111111111110111111111111111111110011111111111111111111111011111111111000111111111111111;
8'h021: data =160'b1111111111111111111000000000000000000000000000000000111111111110011111111111111111011111111111111111111111111111111111111111111111101111111111000111111111111111;
8'h022: data =160'b1111111111111111111100000000000000000000000000000001111111111111111111111111110111111111111111111111111111111111111111111111111111110111111111000111111111111111;
8'h023: data =160'b1111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111000111111111111111;
8'h024: data =160'b1111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111000111111111111111;
8'h025: data =160'b1111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111000111111111111111;
8'h026: data =160'b1111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111000111111111111111;
8'h027: data =160'b1111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111000111111111111111;
8'h028: data =160'b1111111111111111111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111111111111;
8'h029: data =160'b1111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111000111111111111111;
8'h02a: data =160'b1111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111000111111111111111;
8'h02b: data =160'b1111111111111111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111000111111111111111;
8'h02c: data =160'b1111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111000111111111111111;
8'h02d: data =160'b1111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111000111111111111111;
8'h02e: data =160'b1111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110001111000111111111111111;
8'h02f: data =160'b1111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100001111000111111111111111;
8'h030: data =160'b1111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111000001111000111111111111111;
8'h031: data =160'b1111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000011111000111111111111111;
8'h032: data =160'b1111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111000000011111000111111111111111;
8'h033: data =160'b1111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111110000000111111000111111111111111;
8'h034: data =160'b1111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000001111111000111111111111111;
8'h035: data =160'b1111111111111111110001111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111100000000011111111000111111111111111;
8'h036: data =160'b1111111111111110000000001111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111100000000000111111111000111111111111111;
8'h037: data =160'b1111111111111000000001000011111111111111111111000000000000000000000000000001111111111111111111111111111111111111111111100000000000011111111111000111111111111111;
8'h038: data =160'b1111111111110000010001000001111111111111111111110000000000000000000000000000000111111111111111111111111111111111110000000000000001111111111111000111111111111111;
8'h039: data =160'b1111111111100000010001000000111111111111111111111100000000000000000000000000000000000111111111111111111111110000000000000000000111111111111111000111111111111111;
8'h03a: data =160'b1111111111000000011000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000111111111111111;
8'h03b: data =160'b1111111110000000001010100000001111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111000111111111111111;
8'h03c: data =160'b1111111110000000101010100000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000111111111111111;
8'h03d: data =160'b1111111100000000101010100000000111111111111111111111111110000000000001000000000000000000000000000000000000000000000000001111111111111111111111000111111111111111;
8'h03e: data =160'b1111111000000000100010100000000011111111111111111111111111100000000000111000000000000000000000000000000000000000000000011111111111111111111111000111111111111111;
8'h03f: data =160'b1111111000000000100100000000000011111111111111111111111111111000000001001111000000000000000000000000000000000000000000111111111111111111111111000111111111111111;
8'h040: data =160'b1111111000000000000100000000000011111111111111111111111111111000000000010011111000000000000000000000000000000000000001111111111111111111111111000111111111111111;
8'h041: data =160'b1111110000000011000100011000000001111111111111111111111111110000000000001101111111100000000000000000000000000000000011111111111111111111111111000111111111111111;
8'h042: data =160'b1111110000001000000100010110000001111111111111111111111111110000000000000011001111111110000000000000000111000000000111111111111111111111111111000111111111111111;
8'h043: data =160'b1111110000010001000100010001000001111111111111111111111111100010000000111000111001111111111111111111111111000000000011111111111111111111111111000111111111111111;
8'h044: data =160'b1111110000010001000100010001000001111111111111111111111111000111100001111111000111001111111111111111111110000000000001111111111111111111111111000111111111111111;
8'h045: data =160'b1111100000100001000100010000100000111111111111111111111111000111111011111111110000111100111111111111111000000000000000111111111111111111111111000111111111111111;
8'h046: data =160'b1111100000100001000100010000100000111111111111111111111110001111111011111111111110000111111100000000111100000000000000001111111111111111111111000111111111111111;
8'h047: data =160'b1111100000100001000100010000100000111111111111111111111100001111110111111111111111111000000111111111000000000000000000110111111111111111111111000111111111111111;
8'h048: data =160'b1111100000101111000100001100100000111111111111111111111100011111101111111111111111111111111000000000000000000000000000111011111111111111111111000111111111111111;
8'h049: data =160'b1111100000010001000000000011000000111111111111111111111000111111011111111111111111111111111111111000000001100000000000011100111111111111111111000111111111111111;
8'h04a: data =160'b1111100000101000000000000011000000111111111111111111111000111111011111111111111111111111111111111000000111100000000000011111111111111111111111000011111111111111;
8'h04b: data =160'b1111100000100100000010000100100000111111111111111111111001111110111111111111111111111111111111111000111111100000000000011111111110111111011111110110011111111111;
8'h04c: data =160'b1111100001000010001010001000000000111111111111111111111101111101111111111111111111111111111111111011111111100010000000001111111111111110111111111100000111111111;
8'h04d: data =160'b1111100001000001001010010000010000111111111111111111111110111011111111111111111111111111111111111011111111100011000000001111111111111111111111110000000111111111;
8'h04e: data =160'b1111110001000000101010100000010001111111111111111111111111001011111111111111111111111111111111111011111111100011100000000111111111111111111111100000111111111111;
8'h04f: data =160'b1111110000000000101010100000000001111111111111111111111111100111111111111111111111111111111111111011111111100011110000000011111111111111111111000001111111011111;
8'h050: data =160'b1111110000100000010011000000100001111111111111111111111111111111111111111111111111111111111111111011111111100011111000000001111111111101111110000011111111101111;
8'h051: data =160'b1111110000010010001010000001000001111111111111111111111111001111111111111111111111111111111111111011111111110011111100000000011111111100111000000011111111101111;
8'h052: data =160'b1111111000001010001010000010000011111111111111111111111111111000111111111111111111111111111111111011111110000111111110000000001111111100000000000001111111100111;
8'h053: data =160'b1111111000000100001010000000000011111111111111111111111111111111001111111111111111111111111111111000000011101111111111100000000011111100000000000000111111100111;
8'h054: data =160'b1111111100000100001100000100000111111111111111111111111111111111110000011111111111111111111111111111111111111111111111110000000000111000000111100000000011000111;
8'h055: data =160'b1111111100000010001100001000000111111111111111111111111111111111110011100000111111111111111111111111111110001111111111111000000000000000111111111100000000000111;
8'h056: data =160'b1111111110000010000100001000001111111111111111111111111111111111100011111110000000000000111111000000000000101111111111111100000000000001111111111111000000001111;
8'h057: data =160'b1111111110000010000100010000001111111111111111111111111111111111100111111111111110000000000000011111111111110111111111111111000000000001111111111111110000011111;
8'h058: data =160'b1111111111000000000100010000011111111111111111111111111111111111000111111111111111111111111111111111111111111101111111111111100000000000111111111111100001111111;
8'h059: data =160'b1111111111100001000100010000111111111111111111111111111111111111001111111111111001111111111111111111111111111110011111111111111000000000001111111111000001111111;
8'h05a: data =160'b1111111111110001000100010001111111111111111111111111111111111110001111111111111100000011111111111111111111111111101111111111111100000000000000000000000011111111;
8'h05b: data =160'b1111111111111101000100010111111111111111111111111111111111111110011111111111111110000000001111111111111111111111110011111111111111000000000000000000000111111111;
8'h05c: data =160'b1111111111111111000100011111111111111111111111111111111111111100011111111111111111000010000011111111111111111111111101111111111111110000000000000000001111111111;
8'h05d: data =160'b1111111111111111111111111111111111111111111111111111111111111100111111111111111111000011000000111111111111111111111100111111111111111111110000000000011111111111;
8'h05e: data =160'b1111111111111111111111111111111111111111111111111111111111111111000111111111111111000011110000011111111111111111110001111111111111111111111111000111111111111111;
8'h05f: data =160'b1111111111111111111111111111111111111111111111111111111111111111110000001111111111000011111000000111111111111110001110111111111111111111111111000111111111111111;
8'h060: data =160'b1111111111111111111111111111111111111111111111111111111111111111110011110000000000000011111110000001111110000001111111011111111111111111111111000111111111111111;
8'h061: data =160'b1111111111111111111111111111111111111111111111111111111111111111100111111110000000111111111111000000000000011111111111111111111111111111111111000111111111111111;
8'h062: data =160'b1111111111111111111111111111111111111111111111111111111111111111001111111111000000111111111111111110000000011111111111111011111111111111111111000111111111111111;
8'h063: data =160'b1111111111111111111111111111111111111111111111111111111111111111011111111111000000111111111111111111100000001111111111111111111111111111111111000111111111111111;
8'h064: data =160'b1111111111111111111111011111111011111111111111111111111111111110111111111111000000111111111111111111110000000111111111111111011111111111111111000111111111111111;
8'h065: data =160'b1111111111111111011111001101111011111111111111111111111111111110111111111111000000111111111111111111111000000001111111111111110111111111111111000111111111111111;
8'h066: data =160'b1111101111101111111111010111111011111111111111111111111111111101111111111111100000111111111111111111111100000000111111111111111011111111111111110111111111111111;
8'h067: data =160'b1111111111111111111111111111111111111111111111111111111111111001111111111111100000011111111111111111111111000000011111111111111111111111111111111111111111111111;
8'h068: data =160'b1111111111111111111111111111111111111111111111111111111111111011111111111111100000011111111111111111111111100000000111111111111111011111111111111111111111111111;
8'h069: data =160'b1111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111110000000011111111111111110111111111111111111111111111;
8'h06a: data =160'b1111110101111111111110101111011111011111111111111111111111111111111111111110000000111111111111111111111111111000000001111111111111111001111111111111111111111111;
8'h06b: data =160'b1111111101111111111111101011101111111111111111111111111111111111111111111111000000011111111111111111111111111100000000111111111111111111101111111111111111111111;
8'h06c: data =160'b1111111101110111111111101011111101111111111111111111011111111111111111111111000000011111111111111111111111111110000000111111111111111111111100111111111111111111;
8'h06d: data =160'b1111111111111011111111101111111111111111111111111101111111111111111111111111100000011111111111111111111111111111000000011111111111111111111111101111111111111111;
8'h06e: data =160'b1111111111111111111111111111111111111111111111011111111111111100001111111111100000011111111111111111111111111111100000001111111111111111111111111011111111111111;
8'h06f: data =160'b1111111111111111111111111111111111111111111110111111111110000011111111111111000000001111111111111111111111111111110000000111111111111100001111111110111111111111;
8'h070: data =160'b1111111111111111111111111111111111111111111111111111111100011111111111111110000000001111111111111111111111111111111000000001111111111111110011111111110111111111;
8'h071: data =160'b1111101111110111101111011111111111111111111111111111111000111111111111111100000000001111111111111111111111111111111000000000111111111111110001111111111011111111;
8'h072: data =160'b1111111110111111111011011111110111111111111110001111110000111111111111111000000000011111111111111111111111111111111110000000001111111111110001111111111011111111;
8'h073: data =160'b1111101111110111101111011111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111100000001111111111110000111111111011111111;
8'h074: data =160'b1111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111000000000111111100000000000000011111111;
8'h075: data =160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111;
8'h076: data =160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8'h077: data =160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

default : data = 0; 
	endcase
 
 // output logic 
    assign G = data[pix_x_reg[9:2]];
    
endmodule